library verilog;
use verilog.vl_types.all;
entity pratica4 is
    port(
        clock           : in     vl_logic;
        reset           : in     vl_logic
    );
end pratica4;
