module mesi ();

// Instanciar 3 Caches
// Em cada ciclo de clock essas caches serão percorridas


// PASSO A PASSO MESI
// 1) Checar para qual posição da cache a tag indicada está mapeada;
// 2) Se checar se na posição mapeada ocorre read ou write hit ou miss;

endmodule
